

import rfsoc_config::*;


module axis_ps_to_pl
#(parameter ps_axis_width = 32)
(
	input wire clk,
	
	input wire rst,
	
	input wire [15:0] channel_select,
	
	//AXIS input from PS
	input wire [ps_axis_width-1:0] s_axis_tdata,
    input wire s_axis_tvalid,
    output reg s_axis_tready,
	
	
	//AXIS output to PL
	output wire [255:0] m_axis_tdata,
    output wire m_axis_tvalid,
    input wire m_axis_tready
);


parameter ps_per_pl = 256 / ps_axis_width;

reg [15:0] word_cnt;
reg [255:0] word_buff;

//async fifo input bus
reg [255:0] async_fifo_data;
reg async_fifo_valid;
wire async_fifo_ready;



//fifo instantiation
axis_sync_fifo #(4, 256) ps_to_pl_sync_fifo 
(
	rst,
	
	clk,
	async_fifo_valid,
	async_fifo_ready,
	async_fifo_data,

	m_axis_tdata,
	m_axis_tvalid,
	m_axis_tready
	
);

task reset_regs();
begin
	
	async_fifo_data <= 0;
	async_fifo_valid <= 0;
	word_cnt <= 0;
	word_buff <= 0;
	
	s_axis_tready <= 0;

end
endtask

initial begin
	reset_regs();
end

always @ (posedge clk or negedge rst) begin

	if(!rst) begin
	
		reset_regs();
	
	end
	else begin
		
		//Reset write line for async fifo interface
		async_fifo_valid <= 0;
		
		//Always ready to read data till we are not
		s_axis_tready <= 1;

		//if there is an incomming word from PS
		//And a challel is selected
		if(s_axis_tvalid && channel_select != 0) begin
		
			//If this is the last word in the sequence
			if(word_cnt == (ps_per_pl-1)) begin
				//If the async fifo is ready
				if(async_fifo_ready) begin
					//Push this word and the buffer out to the async fifo
					async_fifo_data <= {word_buff[255-ps_axis_width:0], s_axis_tdata};
					word_buff <= {word_buff[255-ps_axis_width:0], s_axis_tdata};
					async_fifo_valid <= 1;
					word_cnt <= 0;
					
					s_axis_tready <= 1;//Indicating we read this word
				end
				else begin
					s_axis_tready <= 0;//Indicating we did not read this word
				end
			end
			else begin
				//Store this word in the correct buffer position
				word_buff <= {word_buff[255-ps_axis_width:0], s_axis_tdata};
				word_cnt <= word_cnt + 1;
			end
		end
		
	end
end




endmodule