

//Routes axis output from PS to one of 16 channels using channel selector